`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:56:56 03/19/2013 
// Design Name: 
// Module Name:    win_checker 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module win_checker(
    input wire [2:0] game_board [0:4][0:4],
    input wire [1:0] player_id,
    output wire player_won,
);

    // TODO: Given player value and game board, determine if that player has won the game
    // player_id = 1 for player 1, 2 for player 2

endmodule